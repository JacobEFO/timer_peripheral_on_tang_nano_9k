/* Copyright (C) reserved for Jacob E. F. Overgaard, 2024
 *
 *
 * @file: timer.v
 * @author: Jacob E. F. Overgaard
 * @date: 2024-07-11
 *
 * @brief:
 *    Timer module that functions as an MCU peripheral
 * 
 */

module uart_rx
(
    input clk_i,
    input rst_ni
);


endmodule //uart_rx
